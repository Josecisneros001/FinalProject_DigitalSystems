library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;

library std;
use std.textio.all;

entity i2c_tb is 
end entity;

architecture arch of i2c_tb is
begin
end arch;