library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_textio.all;

entity i2cTransceiver is
end entity;

architecture arch of i2cTransceiver is
begin
end arch;