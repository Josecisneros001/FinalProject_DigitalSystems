library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity i2cReceiver is 
end entity;

architecture arch of i2cReceiver is
begin
end arch;